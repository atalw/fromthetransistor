// The media-independent interface (MII) is a standard interface to connect a Ethernet media access 
// control (MAC) block to a PHY chip.
// The original MII transfers network data using 4-bit nibbles in each direction (4 transmit data 
// bits, 4 receive data bits). The data is clocked at 25 MHz to achieve 100 Mbit/s throughput.
// https://en.wikipedia.org/wiki/Media-independent_interface
// We're using 8-bit nibbles.
module mii;
    // The transmit clock is a free-running clock generated by the PHY based on the link speed
    // (25 MHz for 100 Mbit/s, 2.5 MHz for 10 Mbit/s).
    // The remaining transmit signals are driven by the MAC synchronously on the rising edge of TXC.
    // This arrangement allows the MAC to operate without having to be aware of the link speed.
    // The transmit enable signal is held high during frame transmission and low when the transmitter
    // is idle.
    wire        w_txc;      // transmit clock
    wire        w_txen;     // transmit enable
    wire [7:0]  w_txd;      // transmit data

    // The first seven receiver signals are entirely analogous to the transmitter signals, except
    // RX_ER is not optional and used to indicate the received signal could not be decoded to valid
    // data. The receive clock is recovered from the incoming signal during frame reception. When
    // no clock can be recovered (i.e. when the medium is silent), the PHY must present a free-running
    // clock as a substitute.
    wire        w_rxc;      // receive clock
    wire        w_rxdv;     // receive data valid
    wire [7:0]  w_rxd;      // receive data
    wire        w_rxer;     // receive error


    mac mac(w_txc, w_rxc, w_rxdv, w_rxd, w_rxer, w_txen, w_txd);

    phy phy(w_txen, w_txd, w_txc, w_rxc, w_rxdv, w_rxd, w_rxer);

endmodule
