module phy_tx(
    input wire in_txen,
    input wire [7:0] in_txd,
    output wire out_txc,
    output wire out_txen,
    output wire [7:0] out_txd
    );

endmodule
