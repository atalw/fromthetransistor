`include "mac.v"
`include "phy.v"

// Encapsulates: Data-link layer <-> MAC <-> MII <-> PHY <-> Wire
// Inputs/Outputs:
// - Higher layer
// - Wire
module eth_controller(
    input   wire          in_txen,      // mcu/cpu to mac transmit enable
    input   wire [7:0]    in_txd,       // mcu/cpu to mac transmit data
    input   wire          in_rxen,      // wire to phy receive enable
    input   wire [7:0]    in_rxd,       // wire to phy receive data
    output  wire          out_tx_ready, // mac to mcu/cpu transmit ready (1 after preamble etc has been sent)
    output  wire          out_dll_rxen, // mac to data-link layer receive enable
    output  wire [7:0]    out_dll_rxd,  // mac to data-link layer receive data
    output  wire          out_wire_txen,// phy to wire transmit enable
    output  wire [7:0]    out_wire_txd  // phy to wire transmit data
    );

    // We've included the MII in this module itself. It is essentially common wires between the MAC
    // and PHY. Since we're instantiating them here, it makes sense to connect them here to.
    //
    // The media-independent interface (MII) is a standard interface to connect a Ethernet media access 
    // control (MAC) block to a PHY chip.
    // The original MII transfers network data using 4-bit nibbles in each direction (4 transmit data 
    // bits, 4 receive data bits). The data is clocked at 25 MHz to achieve 100 Mbit/s throughput.
    // https://en.wikipedia.org/wiki/Media-independent_interface
    //
    // The transmit clock is a free-running clock generated by the PHY based on the link speed
    // (25 MHz for 100 Mbit/s, 2.5 MHz for 10 Mbit/s).
    // The remaining transmit signals are driven by the MAC synchronously on the rising edge of TXC.
    // This arrangement allows the MAC to operate without having to be aware of the link speed.
    // The transmit enable signal is held high during frame transmission and low when the transmitter
    // is idle.
    wire        w_txc;      // transmit clock
    wire        w_txen;     // transmit enable
    wire [7:0]  w_txd;      // transmit data

    // The first seven receiver signals are entirely analogous to the transmitter signals, except
    // RX_ER is not optional and used to indicate the received signal could not be decoded to valid
    // data. The receive clock is recovered from the incoming signal during frame reception. When
    // no clock can be recovered (i.e. when the medium is silent), the PHY must present a free-running
    // clock as a substitute.
    wire        w_rxc;      // receive clock
    wire        w_rxdv;     // receive data valid
    wire [7:0]  w_rxd;      // receive data
    wire        w_rxer;     // receive error
    wire        w_crs;      // carrier sense

    mac mac(
        .in_txc(w_txc),
        .in_txen(in_txen),
        .in_txd(in_txd),
        .in_rxc(w_rxc),
        .in_rxdv(w_rxdv),
        .in_rxd(w_rxd),
        .in_rxer(w_rxer),
        .in_crs(w_crs),
        .out_tx_ready(out_tx_ready),
        .out_txen(w_txen),
        .out_txd(w_txd),
        .out_rxen(out_dll_rxen),
        .out_rxd(out_dll_rxd)
    );

    phy phy(
        .in_txen(w_txen),
        .in_txd(w_txd),
        .in_rxen(in_rxen),
        .in_rxd(in_rxd),
        .out_txc(w_txc),
        .out_txen(out_wire_txen),
        .out_txd(out_wire_txd),
        .out_rxc(w_rxc),
        .out_rxdv(w_rxdv),
        .out_rxd(w_rxd),
        .out_rxer(w_rxer),
        .out_crs(w_crs)
    );

endmodule
